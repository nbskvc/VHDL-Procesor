library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity program_counter is
    Port (
        clk     : in  STD_LOGIC;      
        rst   : in  STD_LOGIC;   
        o_pc  : out STD_LOGIC_VECTOR(15 downto 0);
		  i_pc_clear : in std_logic;
		  i_pc_en : in std_logic
    );
end program_counter;

architecture Behavioral of program_counter is
    signal pc_reg : STD_LOGIC_VECTOR(15 downto 0);
begin

    process(clk, rst)
    begin
        if rst = '0' then
            pc_reg <= (others => '0');  
        elsif rising_edge(clk) then
				if(i_pc_clear = '1')then
					pc_reg <= (others => '0');
				elsif(i_pc_en = '1')then
					if(pc_reg = x"000F")then
						pc_reg <= pc_reg;
					else
						pc_reg <= pc_reg + 1; 
					end if;
				else
					pc_reg <= pc_reg;
				end if;
        end if;
    end process;

    o_pc <= pc_reg;                   

end Behavioral;
